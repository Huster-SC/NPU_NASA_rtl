`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/09/24 11:17:08
// Design Name: 
// Module Name: mac_sim
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mac_sim();
    parameter DATA_WIDTH = 8;
    parameter DATA_NUM   = 32;
     
    reg                                   i_clk      ;
    reg                                   i_rst_n    ;
    reg  [DATA_NUM * DATA_WIDTH-1:0]      i_wdata    ;
    reg                                   i_wdata_vld;
    reg  [DATA_NUM * DATA_WIDTH-1:0]      i_mdata    ;
    reg                                   i_mdata_vld;
    reg                                   i_mac_clear;
    reg                                   i_mac_en;        
    reg  [2:0]                            i_mac_id;
    wire [DATA_NUM * DATA_WIDTH-1:0]      o_wdata    ;
    wire                                  o_wdata_vld;
    wire [DATA_NUM * DATA_WIDTH-1:0]      o_mdata    ;
    wire                                  o_mdata_vld;
    wire [DATA_NUM * 2 * DATA_WIDTH-1:0]  o_mac_result;
    
    wire [5:0] o_count;
    wire [DATA_NUM * DATA_WIDTH - 1:0]  o_r_wdata;
    wire                                o_r_wdata_vld;
    wire [DATA_NUM * DATA_WIDTH - 1:0]  o_r_mdata;
    wire                                o_r_mdata_vld; 
    //input                                               i_mac_clear     ,
    
    pe_mac
    sim_mac(i_clk, i_rst_n, i_mac_en, i_mac_id, i_wdata, i_wdata_vld, i_mdata, i_mdata_vld, i_mac_clear,
            o_wdata, o_wdata_vld, o_mdata, o_mdata_vld, o_mac_result,
            o_count, o_r_wdata, o_r_wdata_vld, o_r_mdata, o_r_mdata_vld);
    
    initial begin 
        i_clk <= 0;
        forever #5 i_clk <= ~i_clk;
    end
    
    initial begin
        i_rst_n  <= 1;
        i_mac_id <= 0;
        i_mac_en <= 1;
    end
    
    initial begin
       i_mdata     <= 0;
       i_mdata_vld <= 0;
       i_wdata     <= 0;
       i_wdata_vld <= 0;
       
       i_mac_clear <= 1;
       #10
       i_mac_clear <= 0;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_mdata_vld <= 1;
       #10
       i_mdata     <= 0;
       i_mdata_vld <= 0;
       
       #20
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201_0201;
       i_wdata_vld <= 1;
       #10
       i_wdata     <= 256'h0;
       i_wdata_vld <= 0;
       
       
    end
    
endmodule
